prac1.cir
.INCLUDE uA741.model
Vcc	4	0	DC	9
Vdd	0	5	DC	9
vg	1	0	DC	0
R1	1	2	10k
R2	2	3	57k
X1	0	2	4	5	3	uA741
.PRINT DC v(3)
.DC vg -2 2 0.1 > grafica.dat
.END
